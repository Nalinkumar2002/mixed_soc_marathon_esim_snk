
module nali_and (a,b,c,d,o);
input a,b,c,d;
output o;

	assign o = a & b & c & d ;

endmodule